module Addcout3 (input [2:0] I0, input [2:0] I1, output [2:0] O, output  COUT);
wire  inst0_O;
wire  inst1_CO;
wire  inst2_O;
wire  inst3_CO;
wire  inst4_O;
wire  inst5_CO;
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst0 (.I0(1'b0), .I1(I0[0]), .I2(I1[0]), .I3(1'b0), .O(inst0_O));
SB_CARRY inst1 (.I0(I0[0]), .I1(I1[0]), .CI(1'b0), .CO(inst1_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst2 (.I0(1'b0), .I1(I0[1]), .I2(I1[1]), .I3(inst1_CO), .O(inst2_O));
SB_CARRY inst3 (.I0(I0[1]), .I1(I1[1]), .CI(inst1_CO), .CO(inst3_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst4 (.I0(1'b0), .I1(I0[2]), .I2(I1[2]), .I3(inst3_CO), .O(inst4_O));
SB_CARRY inst5 (.I0(I0[2]), .I1(I1[2]), .CI(inst3_CO), .CO(inst5_CO));
assign O = {inst4_O,inst2_O,inst0_O};
assign COUT = inst5_CO;
endmodule

module Register3CE (input [2:0] I, output [2:0] O, input  CLK, input  CE);
wire  inst0_Q;
wire  inst1_Q;
wire  inst2_Q;
SB_DFFE inst0 (.C(CLK), .E(CE), .D(I[0]), .Q(inst0_Q));
SB_DFFE inst1 (.C(CLK), .E(CE), .D(I[1]), .Q(inst1_Q));
SB_DFFE inst2 (.C(CLK), .E(CE), .D(I[2]), .Q(inst2_Q));
assign O = {inst2_Q,inst1_Q,inst0_Q};
endmodule

module Counter3CE (output [2:0] O, output  COUT, input  CLK, input  CE);
wire [2:0] inst0_O;
wire  inst0_COUT;
wire [2:0] inst1_O;
Addcout3 inst0 (.I0(inst1_O), .I1({1'b0,1'b0,1'b1}), .O(inst0_O), .COUT(inst0_COUT));
Register3CE inst1 (.I(inst0_O), .O(inst1_O), .CLK(CLK), .CE(CE));
assign O = inst1_O;
assign COUT = inst0_COUT;
endmodule

module Register8CE (input [7:0] I, output [7:0] O, input  CLK, input  CE);
wire  inst0_Q;
wire  inst1_Q;
wire  inst2_Q;
wire  inst3_Q;
wire  inst4_Q;
wire  inst5_Q;
wire  inst6_Q;
wire  inst7_Q;
SB_DFFE inst0 (.C(CLK), .E(CE), .D(I[0]), .Q(inst0_Q));
SB_DFFE inst1 (.C(CLK), .E(CE), .D(I[1]), .Q(inst1_Q));
SB_DFFE inst2 (.C(CLK), .E(CE), .D(I[2]), .Q(inst2_Q));
SB_DFFE inst3 (.C(CLK), .E(CE), .D(I[3]), .Q(inst3_Q));
SB_DFFE inst4 (.C(CLK), .E(CE), .D(I[4]), .Q(inst4_Q));
SB_DFFE inst5 (.C(CLK), .E(CE), .D(I[5]), .Q(inst5_Q));
SB_DFFE inst6 (.C(CLK), .E(CE), .D(I[6]), .Q(inst6_Q));
SB_DFFE inst7 (.C(CLK), .E(CE), .D(I[7]), .Q(inst7_Q));
assign O = {inst7_Q,inst6_Q,inst5_Q,inst4_Q,inst3_Q,inst2_Q,inst1_Q,inst0_Q};
endmodule

module PISO8CE (input  SI, input [7:0] PI, input  LOAD, output  O, input  CLK, input  CE);
wire  inst0_O;
wire  inst1_O;
wire  inst2_O;
wire  inst3_O;
wire  inst4_O;
wire  inst5_O;
wire  inst6_O;
wire  inst7_O;
wire [7:0] inst8_O;
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst0 (.I0(SI), .I1(PI[0]), .I2(LOAD), .I3(1'b0), .O(inst0_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst1 (.I0(inst8_O[0]), .I1(PI[1]), .I2(LOAD), .I3(1'b0), .O(inst1_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst2 (.I0(inst8_O[1]), .I1(PI[2]), .I2(LOAD), .I3(1'b0), .O(inst2_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst3 (.I0(inst8_O[2]), .I1(PI[3]), .I2(LOAD), .I3(1'b0), .O(inst3_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst4 (.I0(inst8_O[3]), .I1(PI[4]), .I2(LOAD), .I3(1'b0), .O(inst4_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst5 (.I0(inst8_O[4]), .I1(PI[5]), .I2(LOAD), .I3(1'b0), .O(inst5_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst6 (.I0(inst8_O[5]), .I1(PI[6]), .I2(LOAD), .I3(1'b0), .O(inst6_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst7 (.I0(inst8_O[6]), .I1(PI[7]), .I2(LOAD), .I3(1'b0), .O(inst7_O));
Register8CE inst8 (.I({inst7_O,inst6_O,inst5_O,inst4_O,inst3_O,inst2_O,inst1_O,inst0_O}), .O(inst8_O), .CLK(CLK), .CE(CE));
assign O = inst8_O[7];
endmodule

module SIPO32CE (input  I, output [31:0] O, input  CLK, input  CE);
wire  inst0_Q;
wire  inst1_Q;
wire  inst2_Q;
wire  inst3_Q;
wire  inst4_Q;
wire  inst5_Q;
wire  inst6_Q;
wire  inst7_Q;
wire  inst8_Q;
wire  inst9_Q;
wire  inst10_Q;
wire  inst11_Q;
wire  inst12_Q;
wire  inst13_Q;
wire  inst14_Q;
wire  inst15_Q;
wire  inst16_Q;
wire  inst17_Q;
wire  inst18_Q;
wire  inst19_Q;
wire  inst20_Q;
wire  inst21_Q;
wire  inst22_Q;
wire  inst23_Q;
wire  inst24_Q;
wire  inst25_Q;
wire  inst26_Q;
wire  inst27_Q;
wire  inst28_Q;
wire  inst29_Q;
wire  inst30_Q;
wire  inst31_Q;
SB_DFFE inst0 (.C(CLK), .E(CE), .D(I), .Q(inst0_Q));
SB_DFFE inst1 (.C(CLK), .E(CE), .D(inst0_Q), .Q(inst1_Q));
SB_DFFE inst2 (.C(CLK), .E(CE), .D(inst1_Q), .Q(inst2_Q));
SB_DFFE inst3 (.C(CLK), .E(CE), .D(inst2_Q), .Q(inst3_Q));
SB_DFFE inst4 (.C(CLK), .E(CE), .D(inst3_Q), .Q(inst4_Q));
SB_DFFE inst5 (.C(CLK), .E(CE), .D(inst4_Q), .Q(inst5_Q));
SB_DFFE inst6 (.C(CLK), .E(CE), .D(inst5_Q), .Q(inst6_Q));
SB_DFFE inst7 (.C(CLK), .E(CE), .D(inst6_Q), .Q(inst7_Q));
SB_DFFE inst8 (.C(CLK), .E(CE), .D(inst7_Q), .Q(inst8_Q));
SB_DFFE inst9 (.C(CLK), .E(CE), .D(inst8_Q), .Q(inst9_Q));
SB_DFFE inst10 (.C(CLK), .E(CE), .D(inst9_Q), .Q(inst10_Q));
SB_DFFE inst11 (.C(CLK), .E(CE), .D(inst10_Q), .Q(inst11_Q));
SB_DFFE inst12 (.C(CLK), .E(CE), .D(inst11_Q), .Q(inst12_Q));
SB_DFFE inst13 (.C(CLK), .E(CE), .D(inst12_Q), .Q(inst13_Q));
SB_DFFE inst14 (.C(CLK), .E(CE), .D(inst13_Q), .Q(inst14_Q));
SB_DFFE inst15 (.C(CLK), .E(CE), .D(inst14_Q), .Q(inst15_Q));
SB_DFFE inst16 (.C(CLK), .E(CE), .D(inst15_Q), .Q(inst16_Q));
SB_DFFE inst17 (.C(CLK), .E(CE), .D(inst16_Q), .Q(inst17_Q));
SB_DFFE inst18 (.C(CLK), .E(CE), .D(inst17_Q), .Q(inst18_Q));
SB_DFFE inst19 (.C(CLK), .E(CE), .D(inst18_Q), .Q(inst19_Q));
SB_DFFE inst20 (.C(CLK), .E(CE), .D(inst19_Q), .Q(inst20_Q));
SB_DFFE inst21 (.C(CLK), .E(CE), .D(inst20_Q), .Q(inst21_Q));
SB_DFFE inst22 (.C(CLK), .E(CE), .D(inst21_Q), .Q(inst22_Q));
SB_DFFE inst23 (.C(CLK), .E(CE), .D(inst22_Q), .Q(inst23_Q));
SB_DFFE inst24 (.C(CLK), .E(CE), .D(inst23_Q), .Q(inst24_Q));
SB_DFFE inst25 (.C(CLK), .E(CE), .D(inst24_Q), .Q(inst25_Q));
SB_DFFE inst26 (.C(CLK), .E(CE), .D(inst25_Q), .Q(inst26_Q));
SB_DFFE inst27 (.C(CLK), .E(CE), .D(inst26_Q), .Q(inst27_Q));
SB_DFFE inst28 (.C(CLK), .E(CE), .D(inst27_Q), .Q(inst28_Q));
SB_DFFE inst29 (.C(CLK), .E(CE), .D(inst28_Q), .Q(inst29_Q));
SB_DFFE inst30 (.C(CLK), .E(CE), .D(inst29_Q), .Q(inst30_Q));
SB_DFFE inst31 (.C(CLK), .E(CE), .D(inst30_Q), .Q(inst31_Q));
assign O = {inst31_Q,inst30_Q,inst29_Q,inst28_Q,inst27_Q,inst26_Q,inst25_Q,inst24_Q,inst23_Q,inst22_Q,inst21_Q,inst20_Q,inst19_Q,inst18_Q,inst17_Q,inst16_Q,inst15_Q,inst14_Q,inst13_Q,inst12_Q,inst11_Q,inst10_Q,inst9_Q,inst8_Q,inst7_Q,inst6_Q,inst5_Q,inst4_Q,inst3_Q,inst2_Q,inst1_Q,inst0_Q};
endmodule

module main (output  D2, output  D1, input  CLKIN, output  TX, input  RX);
wire [7:0] inst0_REC_BYTE;
wire  inst0_TX;
wire  inst0_RECEIVED;
wire [2:0] inst1_O;
wire  inst1_COUT;
wire  inst2_Q;
wire  inst3_O;
wire  inst4_O;
wire  inst5_O;
wire [31:0] inst6_O;
wire  inst7_O;
wire  inst8_CO;
wire  inst9_O;
wire  inst10_CO;
wire  inst11_O;
wire  inst12_CO;
wire  inst13_O;
wire  inst14_CO;
wire  inst15_O;
wire  inst16_CO;
wire  inst17_O;
wire  inst18_CO;
wire  inst19_O;
wire  inst20_CO;
wire  inst21_O;
wire  inst22_CO;
wire  inst23_TX;
receiver inst0 (.iCE_CLK(CLKIN), .RX(RX), .REC_BYTE(inst0_REC_BYTE), .TX(inst0_TX), .RECEIVED(inst0_RECEIVED));
Counter3CE inst1 (.O(inst1_O), .COUT(inst1_COUT), .CLK(CLKIN), .CE(inst4_O));
SB_DFFE inst2 (.C(CLKIN), .E(inst0_RECEIVED), .D(1'b1), .Q(inst2_Q));
SB_LUT4 #(.LUT_INIT(16'h2222)) inst3 (.I0(inst2_Q), .I1(inst1_COUT), .I2(1'b0), .I3(1'b0), .O(inst3_O));
SB_LUT4 #(.LUT_INIT(16'hEEEE)) inst4 (.I0(inst3_O), .I1(inst0_RECEIVED), .I2(1'b0), .I3(1'b0), .O(inst4_O));
PISO8CE inst5 (.SI(1'b1), .PI(inst0_REC_BYTE), .LOAD(1'b1), .O(inst5_O), .CLK(CLKIN), .CE(inst4_O));
SIPO32CE inst6 (.I(inst5_O), .O(inst6_O), .CLK(CLKIN), .CE(inst4_O));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst7 (.I0(1'b0), .I1(inst6_O[8]), .I2(inst6_O[0]), .I3(1'b0), .O(inst7_O));
SB_CARRY inst8 (.I0(inst6_O[8]), .I1(inst6_O[0]), .CI(1'b0), .CO(inst8_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst9 (.I0(1'b0), .I1(inst6_O[9]), .I2(inst6_O[1]), .I3(inst8_CO), .O(inst9_O));
SB_CARRY inst10 (.I0(inst6_O[9]), .I1(inst6_O[1]), .CI(inst8_CO), .CO(inst10_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst11 (.I0(1'b0), .I1(inst6_O[10]), .I2(inst6_O[2]), .I3(inst10_CO), .O(inst11_O));
SB_CARRY inst12 (.I0(inst6_O[10]), .I1(inst6_O[2]), .CI(inst10_CO), .CO(inst12_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst13 (.I0(1'b0), .I1(inst6_O[11]), .I2(inst6_O[3]), .I3(inst12_CO), .O(inst13_O));
SB_CARRY inst14 (.I0(inst6_O[11]), .I1(inst6_O[3]), .CI(inst12_CO), .CO(inst14_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst15 (.I0(1'b0), .I1(inst6_O[12]), .I2(inst6_O[4]), .I3(inst14_CO), .O(inst15_O));
SB_CARRY inst16 (.I0(inst6_O[12]), .I1(inst6_O[4]), .CI(inst14_CO), .CO(inst16_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst17 (.I0(1'b0), .I1(inst6_O[13]), .I2(inst6_O[5]), .I3(inst16_CO), .O(inst17_O));
SB_CARRY inst18 (.I0(inst6_O[13]), .I1(inst6_O[5]), .CI(inst16_CO), .CO(inst18_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst19 (.I0(1'b0), .I1(inst6_O[14]), .I2(inst6_O[6]), .I3(inst18_CO), .O(inst19_O));
SB_CARRY inst20 (.I0(inst6_O[14]), .I1(inst6_O[6]), .CI(inst18_CO), .CO(inst20_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst21 (.I0(1'b0), .I1(inst6_O[15]), .I2(inst6_O[7]), .I3(inst20_CO), .O(inst21_O));
SB_CARRY inst22 (.I0(inst6_O[15]), .I1(inst6_O[7]), .CI(inst20_CO), .CO(inst22_CO));
transmit inst23 (.iCE_CLK(CLKIN), .RX(RX), .transmit_byte({inst21_O,inst19_O,inst17_O,inst15_O,inst13_O,inst11_O,inst9_O,inst7_O}), .TX(inst23_TX));
assign D2 = inst6_O[1];
assign D1 = inst6_O[0];
assign TX = inst23_TX;
endmodule

