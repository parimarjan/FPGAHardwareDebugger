module test(
  input input_byte,
	);

  reg register;

endmodule

  // never resets it.
